** Profile: "SCHEMATIC1-high pass"  [ C:\USERS\SANDIPAN CHAKRABORTY\GOOGLE DRIVE\AIC_Lab\AIC Expt 3-PSpiceFiles\SCHEMATIC1\high pass.sim ] 

** Creating circuit file "high pass.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1 100 1Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
