** Profile: "SCHEMATIC1-qqw"  [ C:\USERS\SANDIPAN CHAKRABORTY\GOOGLE DRIVE\AIC_Lab\AIC-Exp-5-PSpiceFiles\SCHEMATIC1\qqw.sim ] 

** Creating circuit file "qqw.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10m 1m 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
