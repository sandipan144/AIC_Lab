** Profile: "SCHEMATIC1-er"  [ C:\USERS\SANDIPAN CHAKRABORTY\GOOGLE DRIVE\AIC_Lab\WeinsBridge-PSpiceFiles\SCHEMATIC1\er.sim ] 

** Creating circuit file "er.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 30ms 5ms 0.0001 SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
